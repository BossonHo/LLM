module booth_4_multiplier (
    input [7:0] A,        // 8-bit multiplicand (signed)
    input [7:0] B,        // 8-bit multiplier (signed)
    output reg [15:0] P    // 16-bit product
);

    // ... (omitted for brevity) ...