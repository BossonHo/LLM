module parallel_to_serial (
    input wire clk,
    input wire rst,
    input wire [3:0] data_in,
    input wire valid_in,
    output reg serial_out,
    output reg valid_out
);

    reg [3:0] data_buffer;
    reg [2:0] count;

    always @(posedge clk or posedge rst) begin
        if (rst) begin
            data_buffer <= 4'b0;
            count <= 3'b0;
            serial_out <= 1'b0;
            valid_out <= 1'b0;
        end else if (valid_in) begin
            if (count == 3'b0) begin
                data_buffer <= data_in;
                valid_out <= 1'b1;
            end else begin
                serial_out <= data_buffer[3];
                data_buffer <= {data_buffer[2:0], 1'b0};
                count <= count + 1;

                if (count == 4) begin
                    count <= 3'b0;
                    valid_out <= 1'b0;
                end
            end
        end else begin
            valid_out <= 1'b0;
        end
    end

endmodule